module viterbi_top(input clk, input reset, input clk_enable, input [31:0] encoded, output [15:0] Out);
// configuration (3, [6 7])

  Viterbi_Decoder1 u_bit15 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[31]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[30]),  // boolean
                                       .decoded(Out[15])
                                       );
  Viterbi_Decoder1 u_bit14 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[29]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[28]),  // boolean
                                       .decoded(Out[14])
                                       );
  Viterbi_Decoder1 u_bit13 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[27]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[26]),  // boolean
                                       .decoded(Out[13])
                                       );
  Viterbi_Decoder1 u_bit12 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[25]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[24]),  // boolean
                                       .decoded(Out[12])
                                       );
  Viterbi_Decoder1 u_bit11 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[23]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[22]),  // boolean
                                       .decoded(Out[11])
                                       );
  Viterbi_Decoder1 u_bit10 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[21]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[20]),  // boolean
                                       .decoded(Out[10])
                                       );
  Viterbi_Decoder1 u_bit9 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[19]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[18]),  // boolean
                                       .decoded(Out[9])
                                       );
  Viterbi_Decoder1 u_bit8 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[17]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[16]),  // boolean
                                       .decoded(Out[8])
                                       );
  Viterbi_Decoder1 u_bit7 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[15]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[14]),  // boolean
                                       .decoded(Out[7])
                                       );
  Viterbi_Decoder1 u_bit6 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[13]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[12]),  // boolean
                                       .decoded(Out[6])
                                       );
  Viterbi_Decoder1 u_bit5 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[11]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[10]),  // boolean
                                       .decoded(Out[5])
                                       );
  Viterbi_Decoder1 u_bit4 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[9]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[8]),  // boolean
                                       .decoded(Out[4])
                                       );
  Viterbi_Decoder1 u_bit3 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[7]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[6]),  // boolean
                                       .decoded(Out[3])
                                       );
  Viterbi_Decoder1 u_bit2 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[5]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[4]),  // boolean
                                       .decoded(Out[2])
                                       );
  Viterbi_Decoder1 u_bit1 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[3]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[2]),  // boolean
                                       .decoded(Out[1])
                                       );
  Viterbi_Decoder1 u_bit0 (.clk(clk),
                                       .reset(reset),
                                       .enb(clk_enable),
                                       .Viterbi_Decoder1_in_0(encoded[1]),  // boolean
                                       .Viterbi_Decoder1_in_1(encoded[0]),  // boolean
                                       .decoded(Out[0])
                                       );



















endmodule
